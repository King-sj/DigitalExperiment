module tabletFillingMachine(
  input clk
);
endmodule